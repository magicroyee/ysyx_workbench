`timescale 1ns / 1ps
module top(
    
);

    keyboard_sim u_keyboard_sim (
    );

endmodule
