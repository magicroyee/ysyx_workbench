module top(
    
);

    ps2_keyboard u_ps2_keyboard ();

endmodule
